`timescale 1ns/1ps

module or_gate_tb;

reg  a;
reg b;
wire y;

//initiating -- thats what she said
or_gate uut (
    .a(a),
    .b(b),
    .y(y)
);

initial begin 
    $dumpfile("ipor2.vcd");
    $dumpvars(0, or_gate_tb);
    $monitor("%0t | a=%b b=%b | y=%b" , $time, a, b, y);

    //testing -- thats what she did
    a=0; b=0; #10;
    a=0; b=1; #10;
    a=1; b=0; #10;
    a=1; b=1; #10;

    $finish;
end
endmodule